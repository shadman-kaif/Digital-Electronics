* FILE: lab3_l1.sp

********************** begin header *****************************

* Sample Header file for Generic 2.5V 0.25 um process (g25)

.OPTIONS post ACCT OPTS lvltim=2
.OPTIONS post_version=9007

**################################################
* Only Typical/Typical models included
* NEED TO CHANGE ${MMI_TOOLS} TO BE PHYSICAL PATH
.include '/cad2/mmi_local/sue/g25.mod'
* NOTE: these are contrived spice models
**################################################

.param  arean(w,sdd) = '(w*sdd*1p)'
.param  areap(w,sdd) = '(w*sdd*1p)'
* Setup either one or the other of the following
* For ACM=0,2,10,12 fet models
.param  perin(w,sdd) = '(2u*(w+sdd))'
.param  perip(w,sdd) = '(2u*(w+sdd))'
* For ACM=3,13 fet models
*.param  perin(w,sdd) = '(1u*(w+2*sdd))'
*.param  perip(w,sdd) = '(1u*(w+2*sdd))'

.param ln_min   =  0.25u
.param lp_min   =  0.25u

* used in source/drain area/perimeter calculation
.param sdd        =  0.95

.PARAM vddp=2.5		$ VDD voltage

VDD vdd 0 DC vddp 

.TEMP 105
.TRAN 10p 16n
*********************** end header ******************************

* SPICE netlist for "lab3_l1" generated by MMI_SUE5.6.29 on Thu Mar 16 
*+ 14:07:16 EDT 2023.

* start main CELL lab3_l1
* .SUBCKT lab3_l1 Vi Vo 
C_1 GND Vo 0.3pF 
VVdd net_1 GND DC 2.5V 
M_1 Vo Vi net_1 vdd p W='1.5*1u' L=lp_min ad='areap(1.5,sdd)' 
+ as='areap(1.5,sdd)' pd='perip(1.5,sdd)' ps='perip(1.5,sdd)' 
M_2 Vo Vi GND gnd n W='0.5*1u' L=ln_min ad='arean(0.5,sdd)' 
+ as='arean(0.5,sdd)' pd='perin(0.5,sdd)' ps='perin(0.5,sdd)' 
V_1 Vi GND pulse 0 vddp 0ns 200ps 200ps 6ns 12ns 
* .ENDS	$ lab3_l1

.GLOBAL gnd

.END

