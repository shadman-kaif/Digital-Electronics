magic
tech scmos
use /nfs/ug/homes-4/k/kaifmd/mmi_private/tutorial/sue/FA.lvs /nfs/ug/homes-4/k/kaifmd/mmi_private/tutorial/sue/FA.lvs_0
transform 1 0 0 0 1 0
box 0 0 10 10
<< end >>
